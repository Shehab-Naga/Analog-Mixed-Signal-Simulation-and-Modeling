OverDamped RLC Circuit

Vac 1 0 AC 1
R1 1 2 200
L1 2 3 10u
C1 3 0 10n
.AC DEC 10 1 100meg
.END


